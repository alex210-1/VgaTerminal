--! FontTable.vhd
--! Alexander Horstkötter 13.11.2022

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants.all;

entity FontTable is
    port (
        clk, nrst, en : in std_logic;
        char_addr     : in integer range 0 to 255;
        char_x        : in integer range 0 to CHAR_WIDTH - 1;
        char_y        : in integer range 0 to CHAR_HEIGHT - 1;
        pixel         : out std_logic);
end entity;

architecture xilinx7 of FontTable is
    subtype CharType is std_logic_vector(0 to CHAR_SIZE - 1);
    type FontTableArray is array(0 to (256) * CHAR_SIZE - 1) of std_logic;
    type InputBlobArray is array(0 to (256) - 1) of std_logic_vector(0 to CHAR_SIZE - 1);

    -- ye big old blob o' data (fits in 3 BRAMS)
    -- TODO choose better codepage
    constant INPUT_BLOB : InputBlobArray := (
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000000000000000000000006001F803FE0FFF3FFF3FFF3CF930F800F800F800000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000001800180018001800180018001800180018000000000018003C00180000000000000000000000000",
        x"0000000000000E700E700660066006600000000000000000000000000000000000000000000000000000000000000000",
        x"00000000000000000618061806183FFE04300C300C300C300C307FFC1860186018601860000000000000000000000000",
        x"01800180018001800FF81D9C198019801D800F8003F001F8019C018C018C119C3DF80FE0018001800180000000000000",
        x"00000000000000003E06770C6318E33063603EC0018003FC03E606C60CC718C630EE603C000000000000000000000000",
        x"000000000000000007C01C70380038001C0007FE1C18301830187018301830181C700FE0000000000000000000000000",
        x"000000000000018001800180018001800000000000000000000000000000000000000000000000000000000000000000",
        x"00000000006001C00380070006000C000C001C001C001C001C000C000C000E0006000300018000E00020000000000000",
        x"000000000600038001C000E00060003000300038003800380038003000300070006000C0018007000400000000000000",
        x"000000000000000000000000018001800180399C7FFE03C007E00E701C38081000000000000000000000000000000000",
        x"000000000000000000000000018001800180018001803FFC018001800180018000000000000000000000000000000000",
        x"00000000000000000000000000000000000000000000000000000000000003C003C003C0018003800300070000000000",
        x"000000000000000000000000000000000000000000001FF8000000000000000000000000000000000000000000000000",
        x"00000000000000000000000000000000000000000000000000000000000003C003C003C0000000000000000000000000",
        x"000000000006000C001C001800300070006000C001C001800300070006000C001C001800300070000000000000000000",
        x"000000000000000007E00E701C381838385C30CC308C310C330C3A1C1C181C180E7007E0000000000000000000000000",
        x"000000000000000001C007C01EC010C000C000C000C000C000C000C000C000C000C01FFC000000000000000000000000",
        x"00000000000000000FC03CF030300038003800300070006001C0038006000C0038003FF8000000000000000000000000",
        x"00000000000000000FC03CF010380018003800700380007000180018001820387CF00FC0000000000000000000000000",
        x"000000000000010001800300030006000E000C301C30183038303FFC0030003000300030000000000000000000000000",
        x"00000000000000001FF818001800180018001FE01C780018001C001C001810183C700FC0000000000000000000000000",
        x"000000000000000003F80F300C001800180033F03638381C300C380C180C18180E7807E0000000000000000000000000",
        x"00000000000000001FF80018001800300070006000E000C0018001800300070006000E00000000000000000000000000",
        x"000000000000000007E01E781818381C18181C3007E00CF0381C300C300C381C1E7807E0000000000000000000000000",
        x"000000000000000007E01E7038383018301C301C301C1C7C0FD800180038007001E01F80080000000000000000000000",
        x"000000000000000000000000000003C003C003C00000000000000000000003C003C003C0000000000000000000000000",
        x"000000000000000000000000000003C003C003C0000000000000000003C003C003C00180038003000700000000000000",
        x"0000000000000000000000000008003C00F003C00E0038003C000F0003C000F0001C0000000000000000000000000000",
        x"0000000000000000000000000000000000001FF80000000000001FF80000000000000000000000000000000000000000",
        x"00000000000000000000000010003C000F0003C00070001C003C00F003C00F0038000000000000000000000000000000",
        x"000000000000000007E03E7810180018003800F001C00380030000000000038003800380000000000000000000000000",
        x"00000000000000000FE07C78E01C000E00061F8639C670C760C760C760C760C660C671463E46003C0000000000000000",
        x"000000000000000003C003C007E0066006600C300C30183818183FFC300C300C600E6006000000000000000000000000",
        x"00000000000000001FE018781818181C181818381FC01838180C180C180C181C18781FE0000000000000000000000000",
        x"000000000000000003F80F1E1C00180030003000300030003000300018001C040F1E03F8000000000000000000000000",
        x"00000000000000003FC038F03818380C380C380E380E380E380E380C381C381838F03FC0000000000000000000000000",
        x"00000000000000001FFC1C001C001C001C001C001FF01C001C001C001C001C001C001FFC000000000000000000000000",
        x"00000000000000000FFE0C000C000C000C000C000FF80C000C000C000C000C000C000C00000000000000000000000000",
        x"000000000000000003F00F3C180038003000700070FC700C700C300C300C380C1E3C07F0000000000000000000000000",
        x"0000000000000000381C381C381C381C381C381C3FFC381C381C381C381C381C381C381C000000000000000000000000",
        x"00000000000000001FF80180018001800180018001800180018001800180018001801FF8000000000000000000000000",
        x"000000000000000007F8001800180018001800180018001800180018001800383CF00FC0000000000000000000000000",
        x"0000000000000000180E18181830186019C01B801F001B8019C018E018701838181C180F000000000000000000000000",
        x"00000000000000000C000C000C000C000C000C000C000C000C000C000C000C000FFC0FFC000000000000000000000000",
        x"0000000000000000381C3C3C3C3C3C3C3C2C766E666E664E63C663C66386600660066006000000000000000000000000",
        x"00000000000000003C0C3C0C3E0C360C370C330C318C318C30CC30CC306C306C303C303C000000000000000000000000",
        x"000000000000000007E01E78181C300C300C700E700E700E700E300C300C381C1E7807E0000000000000000000000000",
        x"00000000000000001FF0183C180E180E180E180E181C1FF0180018001800180018001800000000000000000000000000",
        x"000000000000000007E01E78181C300C300C700E700E700E700E300C300C38181E7007F0001C000E0007000000000000",
        x"00000000000000001FE01878181C180C180C180C18381FF018C0186018701838181C180E000000000000000000000000",
        x"000000000000000007F01E7C3808300038001E0007E000F8001C000C000C201C7C780FE0000000000000000000000000",
        x"00000000000000007FFE0180018001800180018001800180018001800180018001800180000000000000000000000000",
        x"0000000000000000300C300C300C300C300C300C300C300C300C300C300C38181E7807E0000000000000000000000000",
        x"00000000000000006006700E300C380C181818180C300C300E70066007E003C003C00180000000000000000000000000",
        x"0000000000000000E003E00763C663C663C663C66246366C366C366C366C342C3C381C38000000000000000000000000",
        x"0000000000000000700E18181C380E70066003C0018003C006600E700C301818301C700E000000000000000000000000",
        x"00000000000000007006300C381C1C180C30066007E003C0018001800180018001800180000000000000000000000000",
        x"00000000000000001FFC000C00180030006000E001C00380030006000C00180038003FFC000000000000000000000000",
        x"000007F00600060006000600060006000600060006000600060006000600060006000600060007F00000000000000000",
        x"0000000060003000380018000C000E00060003000380018000C000E00060003000380018000C000E0000000000000000",
        x"00000FE0006000600060006000600060006000600060006000600060006000600060006000600FE00000000000000000",
        x"018003C007E006600C301838381C00000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000007FFE000000000000",
        x"000000000000070003C00060000000000000000000000000000000000000000000000000000000000000000000000000",
        x"00000000000000000000000000000FE01C70003800380FF81C383838303830383CF80F8C000000000000000000000000",
        x"000000000000180018001800180019F01E781C1C181C180C180C180C181C18181E781BE0000000000000000000000000",
        x"000000000000000000000000000003F00F3C1C00180018003800180018001C000F3C03F0000000000000000000000000",
        x"000000000000001800180018001807D81E7818183818301830183018381838181E7807D8000000000000000000000000",
        x"000000000000000000000000000007E00E701818380C300C3FFC3000380018000E3807F0000000000000000000000000",
        x"00000000000000FE03C40300030003003FF8030003000300030003000300030003000300000000000000000000000000",
        x"000000000000000000000000000407FE1C703818301838181C380FE0180018001C000FF8000C300C3C3C0FF000000000",
        x"000000000000180018001800180019F01F381C1818181818181818181818181818181818000000000000000000000000",
        x"00000000010003C00180000000001FC000C000C000C000C000C000C000C000C000C01FFC000000000000000000000000",
        x"00000000004000E00060000000000FF00030003000300030003000300030003000300070006001C00F801C0000000000",
        x"0000000008001800180018001800181C183818E019C01B801F8019C018E018701838180E000000000000000000000000",
        x"0000000000003F00030003000300030003000300030003000300030003000300038800F8000000000000000000000000",
        x"00000000000000000000000000006F3C7BEC718661866186618661866186618661866186000000000000000000000000",
        x"000000000000000000000000000019F01F381C1818181818181818181818181818181818000000000000000000000000",
        x"000000000000000000000000000007E00E781818381C300C300C300C381C18181E7007E0000000000000000000000000",
        x"000000000000000000000000000019F01E781C1C181C180C180C180C181C18181E781BE0180018001800180000000000",
        x"000000000000000000000000000007D81E7818183818301830183018381818181E780FD8001800180018001800000000",
        x"00000000000000000000000000001E7C06EC078C070C0600060006000600060006001FC0000000000000000000000000",
        x"000000000000000000000000000007F01E38180018000F0003F00038001810183C780FE0000000000000000000000000",
        x"00000000000000000300070007003FF007000700070007000700070007000700038801FC000000000000000000000000",
        x"00000000000000000000000000001818181818181818181818181818181818181C780F98000000000000000000000000",
        x"0000000000000000000000000000300C381C181818180C300C300660066003C003C003C0000000000000000000000000",
        x"0000000000000000000000000000E007618663C663C633C6324C366C366C366C14281C38000000000000000000000000",
        x"0000000000000000000000000000381C1C380E70076003C003C003E006600C301818701E000000000000000000000000",
        x"0000000000000000000000000000300C381C181818180C300C3006600660076003C003C00180038007001C0000000000",
        x"00000000000000000000000000001FF800380070006000C00180030006000E001C001FF8000000000000000000000000",
        x"000000F001C001800180018001800180018003801E000380018001800180018001800180018000F00000000000000000",
        x"000001800180018001800180018001800180018001800180018001800180018001800180018001800000000000000000",
        x"00000F00038001800180018001800180018001C0007801C001800180018001800180018001800F000000000000000000",
        x"00000000000000000000000000000000000000001F06338C60F800000000000000000000000000000000000000000000",
        x"000000000000000000007F806180618061806180618061806180618061806180618061807F8000000000000000000000",
        x"000000000000000001FC038C06000C000C007FF01C001C007FE01C000C000E00078C01F8000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000001C003C001C001800380030000000000",
        x"00000000000001F80398030003001FE00300030003000300030003000300030003000300070006000E00180000000000",
        x"00000000000000000000000000000000000000000000000000000000000000000E381E780E380C701C60186000000000",
        x"000000000000000000000000000000000000000000000000000000000000718E73CE718E000000000000000000000000",
        x"00000000000000000180018001803FFC0180018001800180018001800180018001800180000000000000000000000000",
        x"00000000000000000180018001803FFC018001800180018001803FFC0180018001800180000000000000000000000000",
        x"0000000001C007E00C300000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"00000000000000001E007300630063063E7C03C0BC0040003E3C33666343634237661E3C000000000000000000000000",
        x"0C3007E003C0000007F01E7C3808300038001E0007E000F8001C000C000C201C7C780FE0000000000000000000000000",
        x"00000000000000000000000000000000006000C00380070007000300018000C000600000000000000000000000000000",
        x"00000000000000001FFF39C060C0E0E0E060C060C07EC060C060E060E0E060C039801FFF000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"061803F001E000001FFC000C00180030006000E001C00380030006000C00180038003FFC000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"0000000000C001C00180038003C003800000000000000000000000000000000000000000000000000000000000000000",
        x"00000000008003C003C00180038003000300000000000000000000000000000000000000000000000000000000000000",
        x"00000000061806380E301C701E781C700000000000000000000000000000000000000000000000000000000000000000",
        x"0000000004101E781E780E301C7018601840000000000000000000000000000000000000000000000000000000000000",
        x"0000000000000000000000000000000003C007E007E007E003C000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000007FFE000000000000000000000000000000000000000000000000",
        x"00000000000000000000000000000000000000000000FFFF000000000000000000000000000000000000000000000000",
        x"0000000007300DF000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"00000000000000000000FFCE19CA19EA19AA19AA19BA19B2198200000000000000000000000000000000000000000000",
        x"000000000C3007E001C00000000007F01E38180018000F0003F00038001810183C780FE0000000000000000000000000",
        x"000000000000000000000000000000000600030001C000E000E000C00180030006000000000000000000000000000000",
        x"00000000000000000000000000003E3C7766E1C3E1C3C183C1FFC180C1C0E1C073673E3E000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"000000000C3007E001C0000000001FF800380070006000C00180030006000E001C001FF8000000000000000000000000",
        x"00000E700C3000007006300C381C1C180C30066007E003C0018001800180018001800180000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"00000000000000000000000000000000018003C001800000000001800180018001800180018001800180018000000000",
        x"000000000000000000C000C000C007F80E101C0018001800180018001C000E1007F800C000C000C00000000000000000",
        x"000000000000000003F0071C0E000C000C000C003FF00C000C000C000C000C0018003FFC000000000000000000000000",
        x"000000000000000000000000600637EC1E781818381C381C18181C383FFC700E00000000000000000000000000000000",
        x"0000000000000000700E380C18180C300E70066003C01FF8018001801FF8018001800180000000000000000000000000",
        x"000000000180018001800180018001800180000000000000000001800180018001800180018001800000000000000000",
        x"000000000000000003F00E381C001C000F000FE0187818181C180FB003E00030003808301FE000000000000000000000",
        x"0000000000000E700C300000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"0000000007E01C38300C63E666664C024C024C026C066E2637EC1C180FF0000000000000000000000000000000000000",
        x"0000000000000FE008700030003007F01C3018301C700F98000000000000000000001FF8000000000000000000000000",
        x"00000000000000000000000000000000031C06380C7038E038C01CE00E300718030C0000000000000000000000000000",
        x"000000000000000000000000000000000000000000001FF8001800180018000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000FF0000000000000000000000000000000000000000000000000",
        x"00000000000007E01C3837CC2664666667C666C6366C1C380FF000000000000000000000000000000000000000000000",
        x"0000000000000FF000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        x"0000000000001F8039C030C030C038C01F80000000000000000000000000000000000000000000000000000000000000",
        x"00000000000000000000000000000180018001801FF80180018001800180000000001FF8000000000000000000000000",
        x"0000000000000000000007E00E600030006001C006000FF0000000000000000000000000000000000000000000000000",
        x"0000000000000000000007E00C70003001C000300E7007E0000000000000000000000000000000000000000000000000",
        x"00000000002000E007800400000000000000000000000000000000000000000000000000000000000000000000000000",
        x"00000000000000000000000000003818381838183818381838183818381838383CF8379C380038003800380000000000",
        x"00000000000000000FFE3FC63FC67FC67FC63FC63FC607C600C600C600C600C600C600C600C600C600C600C600000000",
        x"000000000000000000000000000000000000000003C003C003C000000000000000000000000000000000000000000000",
        x"000000000000000000000000000000000000000000000000000000000000000000000000018001800060006007C00000",
        x"0000000000000000000000E007E002600060006000600060000000000000000000000000000000000000000000000000",
        x"00000000000007E00C30181818181818181818180C3007E0000000000000000000001FF8000000000000000000000000",
        x"0000000000000000000000000000000038C01C600E30071C031C07380C7018E030C00000000000000000000000000000",
        x"000000000000000018007800D80018001802181E18F003C01E18F030006600C600FF0006000000000000000000000000",
        x"000000000000000018007800D80018001802181E187803C00E3EF8E74003000E0030007F000000000000000000000000",
        x"00000000000000007E00C3001C000300C3077E3801E007183C386030006600C600FF0006000000000000000000000000",
        x"000000000000000000000000000001C001C001C00000000000C000C001C003800E001C001800180C0E7807E000000000",
        x"0200078000E0000003C003C007E0066006600C300C30183818183FFC300C300C600E6006000000000000000000000000",
        x"004001E00700000003C003C007E0066006600C300C30183818183FFC300C300C600E6006000000000000000000000000",
        x"07E00C300000000003C003C007E0066006600C300C30183818183FFC300C300C600E6006000000000000000000000000",
        x"07300DF00000000003C003C007E0066006600C300C30183818183FFC300C300C600E6006000000000000000000000000",
        x"00000E700C30000003C003C007E0066006600C300C30183818183FFC300C300C600E6006000000000000000000000000",
        x"0660066003C0000003C003C007E0066006600C300C30183818183FFC300C300C600E6006000000000000000000000000",
        x"000000000000000007FE0F800D800D80198019C018FE30C030E07FE060606060E070C03F000000000000000000000000",
        x"000000000000000003F80F1E1C00180030003000300030003000300018001C040F1E03F800C000C00030003003E00000",
        x"010003C0007000001FFC1C001C001C001C001C001FF01C001C001C001C001C001C001FFC000000000000000000000000",
        x"002000F0038000001FFC1C001C001C001C001C001FF01C001C001C001C001C001C001FFC000000000000000000000000",
        x"03F00618000000001FFC1C001C001C001C001C001FF01C001C001C001C001C001C001FFC000000000000000000000000",
        x"00000738061800001FFC1C001C001C001C001C001FF01C001C001C001C001C001C001FFC000000000000000000000000",
        x"0200078000E000001FF80180018001800180018001800180018001800180018001801FF8000000000000000000000000",
        x"004001E0070000001FF80180018001800180018001800180018001800180018001801FF8000000000000000000000000",
        x"07E00C30000000001FF80180018001800180018001800180018001800180018001801FF8000000000000000000000000",
        x"00000E700C3000001FF80180018001800180018001800180018001800180018001801FF8000000000000000000000000",
        x"00000000000000003FE038F8381C380C380E380E7F863806380E380E380C381C38F83FC0000000000000000000000000",
        x"07300DF0000000003C0C3C0C3E0C360C370C330C318C318C30CC30CC306C306C303C303C000000000000000000000000",
        x"0200078000E0000007E01E78181C300C300C700E700E700E700E300C300C381C1E7807E0000000000000000000000000",
        x"004001E00700000007E01E78181C300C300C700E700E700E700E300C300C381C1E7807E0000000000000000000000000",
        x"07E00C300000000007E01E78181C300C300C700E700E700E700E300C300C381C1E7807E0000000000000000000000000",
        x"07300DF00000000007E01E78181C300C300C700E700E700E700E300C300C381C1E7807E0000000000000000000000000",
        x"00000E700C30000007E01E78181C300C300C700E700E700E700E300C300C381C1E7807E0000000000000000000000000",
        x"0000000000000000000000000000000000001C38066003C003C006601C38000000000000000000000000000000000000",
        x"000000000038003007F01E78187C304C30CC708E718E718E710E330C320C3E1C1E780FE00C001C000000000000000000",
        x"0200078000E00000300C300C300C300C300C300C300C300C300C300C300C38181E7807E0000000000000000000000000",
        x"004001E007000000300C300C300C300C300C300C300C300C300C300C300C38181E7807E0000000000000000000000000",
        x"07E00C3000000000300C300C300C300C300C300C300C300C300C300C300C38181E7807E0000000000000000000000000",
        x"00000E700C300000300C300C300C300C300C300C300C300C300C300C300C38181E7807E0000000000000000000000000",
        x"004001E0070000007006300C381C1C180C30066007E003C0018001800180018001800180000000000000000000000000",
        x"0000000000000000180018001FF0183C180C180E180E180E180C181C1FF0180018001800000000000000000000000000",
        x"00000000000007E00E7018381830187018C019C018E01878181C180E1806180E199C1BF8000000000000000000000000",
        x"000000000000070003C0006000000FE01C70003800380FF81C383838303830383CF80F8C000000000000000000000000",
        x"00000000002000E00780040000000FE01C70003800380FF81C383838303830383CF80F8C000000000000000000000000",
        x"0000000001C007E00C30000000000FE01C70003800380FF81C383838303830383CF80F8C000000000000000000000000",
        x"0000000007300DF00000000000000FE01C70003800380FF81C383838303830383CF80F8C000000000000000000000000",
        x"0000000000000E700C30000000000FE01C70003800380FF81C383838303830383CF80F8C000000000000000000000000",
        x"000003C00660066003C0000000000FE01C70003800380FF81C383838303830383CF80F8C000000000000000000000000",
        x"00000000000000000000000000007E7C67EE01C301833F8371FFC180C180C1C0E7E73C7E000000000000000000000000",
        x"000000000000000000000000000003F00F3C1C00180018003800180018001C000F3C03F000C000C00030003003E00000",
        x"000000000000070003C00060000007E00E701818380C300C3FFC3000380018000E3807F0000000000000000000000000",
        x"00000000002000E007800400000007E00E701818380C300C3FFC3000380018000E3807F0000000000000000000000000",
        x"0000000001C007E00C300000000007E00E701818380C300C3FFC3000380018000E3807F0000000000000000000000000",
        x"0000000000000E700C300000000007E00E701818380C300C3FFC3000380018000E3807F0000000000000000000000000",
        x"000000000000070003C0006000001FC000C000C000C000C000C000C000C000C000C01FFC000000000000000000000000",
        x"00000000002000E00780040000001FC000C000C000C000C000C000C000C000C000C01FFC000000000000000000000000",
        x"0000000001C007E00C30000000001FC000C000C000C000C000C000C000C000C000C01FFC000000000000000000000000",
        x"0000000000000E700C30000000001FC000C000C000C000C000C000C000C000C000C01FFC000000000000000000000000",
        x"0000000008600FC001C007700630001807DC1C7C381C300C300C300C300C38181E7007E0000000000000000000000000",
        x"0000000007300DF000000000000019F01F381C1818181818181818181818181818181818000000000000000000000000",
        x"000000000000070003C00060000007E00E781818381C300C300C300C381C18181E7007E0000000000000000000000000",
        x"00000000002000E007800400000007E00E781818381C300C300C300C381C18181E7007E0000000000000000000000000",
        x"0000000001C007E00C300000000007E00E781818381C300C300C300C381C18181E7007E0000000000000000000000000",
        x"0000000007300DF000000000000007E00E781818381C300C300C300C381C18181E7007E0000000000000000000000000",
        x"0000000000000E700C300000000007E00E781818381C300C300C300C381C18181E7007E0000000000000000000000000",
        x"000000000000000000000000018003C00180000000001FF800000000018003C001800000000000000000000000000000",
        x"000000000000000000000030003007E00E7018D838DC308C318C310C3B1C1B180E7007E00C000C000000000000000000",
        x"000000000000070003C0006000001818181818181818181818181818181818181C780F98000000000000000000000000",
        x"00000000002000E00780040000001818181818181818181818181818181818181C780F98000000000000000000000000",
        x"0000000001C007E00C30000000001818181818181818181818181818181818181C780F98000000000000000000000000",
        x"0000000000000E700C30000000001818181818181818181818181818181818181C780F98000000000000000000000000",
        x"00000000002000E0078004000000300C381C181818180C300C3006600660076003C003C00180038007001C0000000000",
        x"000000000000180018001800180019F01E781C1C181C180C180C180C181C18181E781BE0180018001800180000000000",
        x"0000000000000E700C3000000000300C381C181818180C300C3006600660076003C003C00180038007001C0000000000"
    );

    function init_ram_from_blob (blob : in InputBlobArray) return FontTableArray is
        variable font                     : FontTableArray;
    begin
        for i_char in blob'range loop
            for i_pixel in 0 to CHAR_SIZE - 1 loop
                font(i_char * CHAR_SIZE + i_pixel) := blob(i_char)(i_pixel);
            end loop;
        end loop;

        return font;
    end function;

    signal FONT_TABLE : FontTableArray := init_ram_from_blob(INPUT_BLOB);
    signal address    : integer range FONT_TABLE'range;
    signal en_delayed : std_logic; --! delay en 1 tick to match address

    -- required to infer block ram, see Xilinx UG901 P.177
    attribute rom_style               : string;
    attribute rom_style of FONT_TABLE : signal is "block";

    -- prevents inference of dsp, which would be overkill und fuck up the timing
    attribute use_dsp            : string;
    attribute use_dsp of xilinx7 : architecture is "no";
begin
    process (clk) begin
        if rising_edge(clk) then
            if nrst = '0' then
                pixel <= '0';
            else
                address    <= char_addr * CHAR_SIZE + char_y * CHAR_WIDTH + char_x;
                en_delayed <= en;

                if en_delayed = '1' then
                    pixel <= FONT_TABLE(address);
                else
                    pixel <= '0';
                end if;
            end if;
        end if;
    end process;
end architecture;